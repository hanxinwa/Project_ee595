`include "uvm_macros.svh"
import uvm_pkg::*;
`include "./SFQ_PKG.sv"
`include "./and_modules.sv"
`include "./buf_modules.sv"
`include "./top_sv.sv"
`include "./interface.sv"
`include "base_driver.sv"
`include "base_sequencer.sv"
`include "base_monitor.sv"