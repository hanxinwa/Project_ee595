`define pw 1

interface and_if;
    SFQ #(`pw) clk();
    SFQ #(`pw) in1();
    SFQ #(`pw) in2();
    SFQ #(`pw) in3();
    SFQ #(`pw) out();
endinterface